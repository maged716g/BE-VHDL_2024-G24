
module Sopc_Cap (
	clk_clk,
	avalon_cap_0_in_pwm_compas_beginbursttransfer);	

	input		clk_clk;
	input		avalon_cap_0_in_pwm_compas_beginbursttransfer;
endmodule
